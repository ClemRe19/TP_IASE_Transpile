module and_gate3 (e1, e2, e3, s);
    input e1;
    input e2;
    input e3;
    output s;


    assign s = e1 & e2 & e3;

endmodule


//module reg_lin(X, s):



//end module