module add_8_bit (e1, e2, s);
    input [7:0] e1, e2;
    
    output [7:0] s; 

    assign s = e1 + e2;

endmodule


//module reg_lin(X, s):



//end module